-- package for defining generic parameters and signal types
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.fixed_pkg.all;
use IEEE.std_logic_signed.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;

package fir_fixed_generics_package is
    constant ORDER              : integer := 50;
    constant BIT_WIDTH          : integer := 16;
    constant AXIS_WIDTH         : integer := 32;
    constant FRACTIONAL_WIDTH   : integer := 15; -- BIT_WIDTH - 1
    constant COEFFICIENT_WIDTH  : integer := 16; 
    constant COEFFICIENT_LENGTH : integer := (integer(floor(real(ORDER/2))) + 1)*COEFFICIENT_WIDTH;
    constant COEFFICIENT_NUMBER : integer := integer(floor(real(ORDER/2)));
    constant FIFO_DELAY         : integer := 1;
    constant PIPE_DELAY         : integer := COEFFICIENT_NUMBER + 4;
    type reg_array is array(natural range <>) of sfixed(BIT_WIDTH-FRACTIONAL_WIDTH-1 downto -FRACTIONAL_WIDTH);
    type coefficient_fixed_array is array(0 to COEFFICIENT_NUMBER) of sfixed(COEFFICIENT_WIDTH-FRACTIONAL_WIDTH-1 downto -FRACTIONAL_WIDTH);
    constant FIXED_COEFFICIENTS  : coefficient_fixed_array := (
        to_sfixed(0.00810390534100997, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(0.0139939370603132, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(0.0189108907005556, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(0.0218035375226890, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(0.0217399615153303, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(0.0180710347968490, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(0.0105770108900642, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(-0.000425370764916858, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(-0.0140346086299292, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(-0.0287881031065154, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(-0.0427623447120998, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(-0.0537444050649743, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(-0.0594596869136981, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(-0.0578323820105221, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(-0.0472491150953144, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(-0.0267937558959265, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(0.00357712978653458, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(0.0429432458347234, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(0.0894300811571629, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(0.140323745741493, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(0.192283467119808, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(0.241632137861872, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(0.284695370994223, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(0.318152911276251, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(0.339363873552125, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        to_sfixed(0.346629513548268, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH)
    );
end package fir_fixed_generics_package;


        -- to_sfixed(-0.00101955892407069046, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(-0.00065255563728391084, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(0.00040432153191682566, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(0.00154680883851784239, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(0.00168035385481241605, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(-0.00000000000000000196, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(-0.00277670657191815681, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(-0.00415446275048169528, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(-0.00169993772383667885, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(0.00402808043882074522, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(0.00845070298371066939, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(0.00607046404166685597, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(-0.00387098195557225274, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(-0.01436517348355667578, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(-0.01467361728483655009, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(0.00000000000000000798, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(0.02107520378572750805, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(0.02978972907394649913, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(0.01171935673280114810, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(-0.02732117678633463886, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(-0.05812427795715576634, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(-0.04415493856538225959, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(0.03175871620101571036, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(0.14931951643540891661, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(0.25682768876447192863, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH),
        -- to_sfixed(0.30028488991522439555, BIT_WIDTH-FRACTIONAL_WIDTH-1, -FRACTIONAL_WIDTH)

        